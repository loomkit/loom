module main

import installer

fn main() {
	mut app := installer.app()

	app.run()
}
