module main

fn main() {
	println('Welcome to Loom !')
}
